//////////////////////////////////////////////////////////////////////////////////
// The Cooper Union
// ECE 251 Spring 2024
// Engineer: Jason Hao and Daniel Park
// 
//     Create Date: 2023-02-07
//     Module Name: tb_alu
//     Description: Test bench for simple behavorial ALU
//
// Revision: 1.0 - Initial build
//
//////////////////////////////////////////////////////////////////////////////////
`ifndef TB_ALU
`define TB_ALU

`timescale 1ns/100ps
`include "alu.sv"

module tb_alu;
    parameter n = 16;

    logic [(n-1):0] a, b, s;
    logic [2:0] op;
    logic Zero;

    initial begin
	$dumpfile("alu.vcd");
        $dumpvars(0, uut);
        $monitor("a = %b b = %b op = %b, s = %b, zero = %b", a, b, op, s, Zero);
    end

    initial begin
        //testing op 000
	a <= 16'b0000000000000000;
	b <= 16'b0000000000000000;
	op <= 3'b000;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0011101001001100;

	#10 a <= 16'b0000000000000000;
	#10 a <= 16'b1101010001011101;
        
	//testing op 001
	#10 a <= 16'b0000000000000000;
	b <= 16'b0000000000000000;
	op <= 3'b001;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0011101001001100;

	#10 a <= 16'b0000000000000000;
	#10 a <= 16'b1101010001011101;

        //testing op 010
	#10 a <= 16'b0000000000000000;
	b <= 16'b0000000000000000;
	op <= 3'b010;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0011101001001100;

	#10 a <= 16'b0000000000000000;
	#10 a <= 16'b1101010001011101;

        //testing op 011
	#10 a <= 16'b0000000000000000;
	b <= 16'b0000000000000000;
	op <= 3'b011;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0011101001001100;

	#10 a <= 16'b0000000000000000;
	#10 a <= 16'b1101010001011101;

	//testing op 100
	#10 a <= 16'b0111111111111111;
	b <= 16'b0110001111001101;
	op <= 3'b100;

	#10 a <= 16'b0000000000011011;
	b <= 16'b1111111111111111;

	#10 a <= 16'b1111111111111111;
	b <= 16'b1010001110010010;

	#10 a <= 16'b1010101010101010;
	b <= 16'b1010101010101010;

	//testing op 101
	#10 a <= 16'b0111111111111111;
	b <= 16'b0110001111001101;
	op <= 3'b101;

	#10 a <= 16'b0000000000011011;
	b <= 16'b1111111111111111;

	#10 a <= 16'b1111111111111111;
	b <= 16'b1010001110010010;

	#10 a <= 16'b0000000000000011;
	b <= 16'b1111111111111101;

	//testing op 110
	#10 a <= 16'b0000000000000011;
	b <= 16'b0000000000000010;
	op <= 3'b110;

	#10 a <= 16'b0011100010100101;
	b <= 16'b0100101010010011;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0000000000000001;

	#10 a <= 16'b0000000010101111;
	b <= 16'b1000100101101010;

	//testing op 111
	#10 a <= 16'b0101010111110011;
	b <= 16'b0000000000000111;
	op <= 3'b111;

	#10 a <= 16'b1111111111111111;
	b <= 16'b0000000000000001;
	
	#10 a <= 16'b0101000010010110;
	b <= 16'b0000000000001001;

	#10 a <= 16'b1010110101110101;
	b <= 16'b0000000000000100;

    end

    alu uut(.srca(a), .srcb(b), .opcode(op), .out(s), .zero(Zero));

endmodule
`endif // TB_ALU
